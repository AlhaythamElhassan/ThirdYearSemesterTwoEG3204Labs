library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity programable_4bits_counter is 
	port (
		);
end programable_4bits_counter;

architecture behavioural of programable_4bits_counter is 
begin

edn behavioural;